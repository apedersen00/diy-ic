** sch_path: /home/andreasp/diy-ic/testbench/folded_cascode_tb.sch
**.subckt folded_cascode_tb
C1 voutm GND 100f m=1
C2 voutp GND 100f m=1
V2 vdd GND DC 3.3
V3 vinm GND DC 1.65 AC -1.0
V4 vinp GND DC 1.65 AC 1.0
L9 voutp vinp 4G m=1
C3 vinp GND 4G m=1
L11 voutm vinm 4G m=1
C4 vinm GND 4G m=1
x1 vdd voutp voutm vinp vinm GND folded_cascode
**** begin user architecture code

.lib cornerMOShv.lib mos_tt



.param temp=27
.include folded_cascode_tb.save

.control
op
save all
print @n.x1.xm1.nsg13_hv_nmos[ids]
write folded_cascode_tb.raw
set appendwrite #writing into the same raw file
ac dec 100 1 10e6
save all
let vout = abs(v(voutp) - v(voutm))
let Av = db(v(voutp))
let phase = 180*cph(vout)/pi
write folded_cascode_tb.raw
.endc


**** end user architecture code
**.ends

* expanding   symbol:  folded_cascode.sym # of pins=6
** sym_path: /home/andreasp/diy-ic/schematic/folded_cascode.sym
** sch_path: /home/andreasp/diy-ic/schematic/folded_cascode.sch
.subckt folded_cascode VDD vop von vip vin VSS
*.ipin VDD
*.ipin vip
*.ipin vin
*.opin vop
*.opin von
*.ipin VSS
XM1 net2 vip net1 net1 sg13_hv_nmos w=44u l=1u ng=10 m=11
XM4 net2 pbias_upper VDD VDD sg13_hv_pmos w=57u l=2u ng=10 m=10
XM2 net3 vin net1 net1 sg13_hv_nmos w=44u l=1u ng=10 m=11
XM3 net1 tail_bias VSS VSS sg13_hv_nmos w=10.5u l=1u ng=10 m=10
XM5 net3 pbias_upper VDD VDD sg13_hv_pmos w=57u l=2u ng=10 m=10
XM6 von pbias_lower net2 net2 sg13_hv_pmos w=15u l=1u ng=5 m=10
XM7 vop pbias_lower net3 net3 sg13_hv_pmos w=15u l=1u ng=5 m=10
XM9 vop nbias_upper net5 net5 sg13_hv_nmos w=38u l=5u ng=5 m=10
XM8 von nbias_upper net4 net4 sg13_hv_nmos w=38u l=5u ng=5 m=10
XM11 net5 nbias_lower VSS VSS sg13_hv_nmos w=38u l=5u ng=5 m=10
XM10 net4 nbias_lower VSS VSS sg13_hv_nmos w=38u l=5u ng=5 m=10
V1 tail_bias VSS 1.00
V2 pbias_upper VSS 2.2
V3 pbias_lower VSS 1.5
V4 nbias_upper VSS 1.8
V5 nbias_lower VSS 0.9
.ends

.GLOBAL GND
.end
